** Profile: "SCHEMATIC1-dswaf"  [ E:\P1_2024_433E_Popescu_Vlad_Gabriel_GSD_22_Simulator\Schematics\sch_sim-pspicefiles\schematic1\dswaf.sim ] 

** Creating circuit file "dswaf.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../lib_modelepspice_anexa_1/modele_a1_lib/bc856b.lib" 
.LIB "../../../lib_modelepspice_anexa_1/modele_a1_lib/bc846b.lib" 
.LIB "../../../lib_modelepspice_anexa_1/modele_a1_lib/bc817-25.lib" 
.LIB "../../../lib_modelepspice_anexa_1/modele_a1_lib/bc807-25.lib" 
.LIB "../../../lib_modelepspice_anexa_1/modele_a1_lib/1n4148.lib" 
* From [PSPICE NETLIST] section of C:\Users\Popescu Gabriel\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.TRAN  0 3m 0 10u 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
